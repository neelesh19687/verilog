`timescale 1ns/1ns
`include "andgate.v"

module andgate_tb (
    
);

    reg a,b;
    wire c;

    
    
endmodule